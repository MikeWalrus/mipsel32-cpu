module axi_crossbar_1x2(
        input aclk,
        input aresetn,
        input [3:0] s_axi_awid,
        input [31:0] s_axi_awaddr,
        input [3:0] s_axi_awlen,
        input [2:0] s_axi_awsize,
        input [1:0] s_axi_awburst,
        input [1:0] s_axi_awlock,
        input [3:0] s_axi_awcache,
        input [2:0] s_axi_awprot,
        input [3:0] s_axi_awqos,
        input [0:0] s_axi_awvalid,
        output [0:0] s_axi_awready,
        input [3:0] s_axi_wid,
        input [31:0] s_axi_wdata,
        input [3:0] s_axi_wstrb,
        input [0:0] s_axi_wlast,
        input [0:0] s_axi_wvalid,
        output [0:0] s_axi_wready,
        output [3:0] s_axi_bid,
        output [1:0] s_axi_bresp,
        output [0:0] s_axi_bvalid,
        input [0:0] s_axi_bready,
        input [3:0] s_axi_arid,
        input [31:0] s_axi_araddr,
        input [3:0] s_axi_arlen,
        input [2:0] s_axi_arsize,
        input [1:0] s_axi_arburst,
        input [1:0] s_axi_arlock,
        input [3:0] s_axi_arcache,
        input [2:0] s_axi_arprot,
        input [3:0] s_axi_arqos,
        input [0:0] s_axi_arvalid,
        output [0:0] s_axi_arready,
        output [3:0] s_axi_rid,
        output [31:0] s_axi_rdata,
        output [1:0] s_axi_rresp,
        output [0:0] s_axi_rlast,
        output [0:0] s_axi_rvalid,
        input [0:0] s_axi_rready,
        output [7:0] m_axi_awid,
        output [63:0] m_axi_awaddr,
        output [7:0] m_axi_awlen,
        output [5:0] m_axi_awsize,
        output [3:0] m_axi_awburst,
        output [3:0] m_axi_awlock,
        output [7:0] m_axi_awcache,
        output [5:0] m_axi_awprot,
        output [7:0] m_axi_awqos,
        output [1:0] m_axi_awvalid,
        input [1:0] m_axi_awready,
        output [7:0] m_axi_wid,
        output [63:0] m_axi_wdata,
        output [7:0] m_axi_wstrb,
        output [1:0] m_axi_wlast,
        output [1:0] m_axi_wvalid,
        input [1:0] m_axi_wready,
        input [7:0] m_axi_bid,
        input [3:0] m_axi_bresp,
        input [1:0] m_axi_bvalid,
        output [1:0] m_axi_bready,
        output [7:0] m_axi_arid,
        output [63:0] m_axi_araddr,
        output [7:0] m_axi_arlen,
        output [5:0] m_axi_arsize,
        output [3:0] m_axi_arburst,
        output [3:0] m_axi_arlock,
        output [7:0] m_axi_arcache,
        output [5:0] m_axi_arprot,
        output [7:0] m_axi_arqos,
        output [1:0] m_axi_arvalid,
        input [1:0] m_axi_arready,
        input [7:0] m_axi_rid,
        input [63:0] m_axi_rdata,
        input [3:0] m_axi_rresp,
        input [1:0] m_axi_rlast,
        input [1:0] m_axi_rvalid,
        output [1:0] m_axi_rready
    );
    wire clk = aclk;
    wire rst = ~aresetn;

    wire [15:0] m_axi4_awlen;
    assign m_axi_awlen[7:4] = m_axi4_awlen[11:8];
    assign m_axi_awlen[3:0] = m_axi4_awlen[3:0];
    wire [15:0] m_axi4_arlen;
    assign m_axi_arlen[7:4] = m_axi4_arlen[11:8];
    assign m_axi_arlen[3:0] = m_axi4_arlen[3:0];

    axi_crossbar #
        (
            .M_COUNT(2),
            .S_COUNT(1),
            .S_ID_WIDTH(4),
            .M_REGIONS(8),
            .M_BASE_ADDR({512'hbfc00000_a0000000_00000000_c0000000_40000000_80000000_20000000_1fc00000_ffffffff_ffffffff_ffffffff_ffffffff_ffffffff_ffffffff_bfaf0000_1faf0000}),
            .M_ADDR_WIDTH({32'd22, 32'd28, 32'd28, 32'd30, 32'd30, 32'd29, 32'd29, 32'd22, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd0, 32'd 16, 32'd16})
        ) axi_crossbar (
            .clk              ( clk     ), // i, 1
            .rst            ( rst   ), // i, 1

            .s_axi_arid(s_axi_arid),
            .s_axi_araddr(s_axi_araddr),
            .s_axi_arlen({4'b0, s_axi_arlen}),
            .s_axi_arsize(s_axi_arsize),
            .s_axi_arburst(s_axi_arburst),
            .s_axi_arlock(1'b0),
            .s_axi_arcache(s_axi_arcache),
            .s_axi_arprot(s_axi_arprot),
            .s_axi_arqos(s_axi_arqos),
            .s_axi_arvalid(s_axi_arvalid),
            .s_axi_arready(s_axi_arready),
            .s_axi_rid(s_axi_rid),
            .s_axi_rdata(s_axi_rdata),
            .s_axi_rresp(s_axi_rresp),
            .s_axi_rlast(s_axi_rlast),
            .s_axi_rvalid(s_axi_rvalid),
            .s_axi_rready(s_axi_rready),
            .s_axi_awid(s_axi_awid),
            .s_axi_awaddr(s_axi_awaddr),
            .s_axi_awlen({4'b0, s_axi_awlen}),
            .s_axi_awsize(s_axi_awsize),
            .s_axi_awburst(s_axi_awburst),
            .s_axi_awlock(0),
            .s_axi_awcache(s_axi_awcache),
            .s_axi_awprot(s_axi_awprot),
            .s_axi_awqos(s_axi_awqos),
            .s_axi_awvalid(s_axi_awvalid),
            .s_axi_awready(s_axi_awready),
            .s_axi_wdata(s_axi_wdata),
            .s_axi_wstrb(s_axi_wstrb),
            .s_axi_wlast(s_axi_wlast),
            .s_axi_wvalid(s_axi_wvalid),
            .s_axi_wready(s_axi_wready),
            .s_axi_bid(s_axi_bid),
            .s_axi_bresp(s_axi_bresp),
            .s_axi_bvalid(s_axi_bvalid),
            .s_axi_bready(s_axi_bready),

            .m_axi_arid(m_axi_arid),
            .m_axi_araddr(m_axi_araddr),
            .m_axi_arlen(m_axi4_arlen),
            .m_axi_arsize(m_axi_arsize),
            .m_axi_arburst(m_axi_arburst),
            .m_axi_arlock(),
            .m_axi_arcache(m_axi_arcache),
            .m_axi_arprot(m_axi_arprot),
            .m_axi_arqos(m_axi_arqos),
            .m_axi_arvalid(m_axi_arvalid),
            .m_axi_arready(m_axi_arready),
            .m_axi_rid(m_axi_rid),
            .m_axi_rdata(m_axi_rdata),
            .m_axi_rresp(m_axi_rresp),
            .m_axi_rlast(m_axi_rlast),
            .m_axi_rvalid(m_axi_rvalid),
            .m_axi_rready(m_axi_rready),
            .m_axi_awid(m_axi_awid),
            .m_axi_awaddr(m_axi_awaddr),
            .m_axi_awlen(m_axi4_awlen),
            .m_axi_awsize(m_axi_awsize),
            .m_axi_awburst(m_axi_awburst),
            .m_axi_awlock(),
            .m_axi_awcache(m_axi_awcache),
            .m_axi_awprot(m_axi_awprot),
            .m_axi_awqos(m_axi_awqos),
            .m_axi_awvalid(m_axi_awvalid),
            .m_axi_awready(m_axi_awready),
            .m_axi_wdata(m_axi_wdata),
            .m_axi_wstrb(m_axi_wstrb),
            .m_axi_wlast(m_axi_wlast),
            .m_axi_wvalid(m_axi_wvalid),
            .m_axi_wready(m_axi_wready),
            .m_axi_bid(m_axi_bid),
            .m_axi_bresp(m_axi_bresp),
            .m_axi_bvalid(m_axi_bvalid),
            .m_axi_bready(m_axi_bready)
        );
endmodule
