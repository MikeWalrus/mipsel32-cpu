`define ENTRY 5'd0
`define ENTRYLO0 5'd2
`define ENTRYLO1 5'd3
`define BADVADDR 5'd8
`define COUNT 5'd9
`define ENTRYHI 5'd10
`define COMPARE 5'd11
`define STATUS 5'd12
`define CAUSE 5'd13
`define EPC 5'd14
`define CONFIG 5'd16
